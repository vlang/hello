module hello

// 1
pub fn sayhi() {
  println('hello world from module "hello"')
}
