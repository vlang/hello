module hello

pub fn sayhi() {
  println('hello world from module "hello"')
}
