module hello

// 2
pub fn sayhi() {
  println('hello world from module "hello"')
}
