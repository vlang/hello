module hello

fn sayhi() {
  println('hello world from module hello')
}
