module hello

// 4
pub fn sayhi() {
  println('hello world from module "hello"')
}
