module hello

// 3
pub fn sayhi() {
  println('hello world from module "hello"')
}
